// Copyright (C) 2021  Antmicro
// SPDX-License-Identifier: Apache-2.0
module constants (output out0, output out1);
    assign out0 = 1'b0;
    assign out1 = 1'b1;
endmodule
