module simple_core_2 (
    input wire a,
    output wire y,
    output wire c
);

endmodule
