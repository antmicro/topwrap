module simple_core_1 (
    input wire clk,
    input wire rst,
    output reg z
);

endmodule
